module datapath(clk, rst, regdst, jump, branch, memread, memtoreg, aluop, memwrite, alusrc, regwrite)
    
endmodule