module aluctrltest();
    
endmodule